----------------------------------------------------------------------------------
-- Company: Ruder Boskovic Institute
-- Engineer: Ivan Sovic
-- 
-- Create Date:    02:47:29 08/10/2014 
-- Design Name: 
-- Module Name:    memcontroler - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: A controller device which takes 4 input values of the decomposed image, performs decimation,
-- compression and storing to the output RAM. Implements a state machine. Decimation is controled by signals
-- generated by the Control Unit. Compression is performed by thresholding the decomposed pixel values, and
-- counting the pixels under the threshold. LL component of the image is not compressed but stored raw, while
-- LH, HL and HH components are encoded by two byte values: number of pixels under the threshold, followed by
-- the value of the pixel that follows the count of invalid pixels. A special case is when the count of invalid
-- pixels exceeds 255, then the first value equals 255, and the following value is equal to 0 (this is required
-- to avoid overflow).

--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity memcontroler is
	Generic	(	THRESHOLD : integer := 10;
					DATA_WIDTH : integer := 8;
					ADDR_WIDTH : integer := 16;
					IMAGE_WIDTH : integer := 256;
					IMAGE_HEIGHT : integer := 256
				);
	Port	(	
				clk : in STD_LOGIC;
				en : in STD_LOGIC;
				reset : in  STD_LOGIC;
				
				inLL : in STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				inLH : in STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				inHL : in STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				inHH : in STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				
				rowReady : in STD_LOGIC;
				columnReady : in STD_LOGIC;
				
				address : out STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0);
				dataOut : out STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				dataIn : in STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);
				weOut : out STD_LOGIC;
				
				compressedDataSize : out STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0);
				
				cuFinishedProcessing : in STD_LOGIC;
				finishedCompressing : out STD_LOGIC;
				
				readyForNextData : out STD_LOGIC
			);
end memcontroler;

architecture Behavioral of memcontroler is
	type states is (	stateReset,
							stateWaitForRowAndColumn,
							stateProcessData,
							
							stateProcessLL, stateProcessLLIncreaseSP,
							
							stateProcessLH, stateProcessLHCount,
							stateProcessLHSend1, stateProcessLHIncreaseSP1,
							stateProcessLHSend2, stateProcessLHIncreaseSP2, stateProcessLHClearCount,

							stateProcessHL, stateProcessHLCount, stateProcessHLSend1, stateProcessHLIncreaseSP1,
							stateProcessHLSend2, stateProcessHLIncreaseSP2, stateProcessHLClearCount,

							stateProcessHH, stateProcessHHCount, stateProcessHHSend1, stateProcessHHIncreaseSP1,
							stateProcessHHSend2, stateProcessHHIncreaseSP2, stateProcessHHClearCount,
							
							stateSendRemainingData,
							stateSendRemainingDataLH1, stateSendRemainingDataLHIncreaseSP1,
							stateSendRemainingDataLH2, stateSendRemainingDataLHIncreaseSP2,
							stateSendRemainingDataLHClearCount,
							
							stateSendRemainingDataHL1, stateSendRemainingDataHLIncreaseSP1,
							stateSendRemainingDataHL2, stateSendRemainingDataHLIncreaseSP2,
							stateSendRemainingDataHLClearCount,

							stateSendRemainingDataHH1, stateSendRemainingDataHHIncreaseSP1,
							stateSendRemainingDataHH2, stateSendRemainingDataHHIncreaseSP2,
							stateSendRemainingDataHHClearCount,
							
							stateMoveHL, stateMoveHLCheckDone, stateMoveHLSetAddressRead, stateMoveHLReadData, stateMoveHLIncreaseSP,
							stateMoveHH, stateMoveHHCheckDone, stateMoveHHSetAddressRead, stateMoveHHReadData, stateMoveHHIncreaseSP,
							
							stateSendData, stateSendData2,
							stateFinished, stateFinished2, stateFinished3);

	signal currentState : states := stateReset;
	signal nextState : states := stateReset;
	signal returnState : states := stateReset;
	
	constant totalNumPixels : integer := IMAGE_WIDTH * IMAGE_HEIGHT;
	constant spLLTop : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := (others => '0');
	constant spLHTop : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := conv_std_logic_vector((1*(totalNumPixels /4)), ADDR_WIDTH);
	constant spHLTop : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := conv_std_logic_vector((2*(totalNumPixels /4)), ADDR_WIDTH);
	constant spHHTop : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := conv_std_logic_vector((3*(totalNumPixels /4)), ADDR_WIDTH);
	
	-- Stack pointer initialization
	signal spLL : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spLLTop;
	signal spLH : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spLHTop;
	signal spHL : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spHLTop;
	signal spHH : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spHHTop;
	
	signal spHLMoving : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spHLTop;
	signal spHHMoving : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := spHHTop;
	
	signal sameCountLH : integer := 0;
	signal sameCountHL : integer := 0;
	signal sameCountHH : integer := 0;
	
	signal dataToSend : STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0) := (others => '0');
	signal addressToSend : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) downto 0) := (others => '0');
	signal receivedData : STD_LOGIC_VECTOR((DATA_WIDTH - 1) downto 0);

begin
	process (clk, reset, nextState)
	begin
		if reset = '1' then
			currentState <= stateReset;
		elsif rising_edge(clk) then
			if en = '1' then
				-- Perform all synchronous signal changes. These are changes that
				-- cannot be performed in the combinational process because they
				-- would infer the usage of implicit latches. Example of such a signal
				-- is spLL which counts the current address of the data to be stored
				-- (stack pointer).
				if currentState <= stateReset then								-- Initialize all stack pointers and counters.
					spLL <= spLLTop;
					spLH <= spLHTop;
					spHL <= spHLTop;
					spHH <= spHHTop;
					sameCountLH <= 0;
					sameCountHL <= 0;
					sameCountHH <= 0;
					
				
				-----------------------------------------------------------------
				-- These states are used for counting the values that are
				-- lower than the given threshold, and storing the results
				-- to the output RAM. These states occur while
				-- cuFinishedProcessing is low.
				-----------------------------------------------------------------
				-----
				-- Process the LL component of the image. This consists simply of storing the raw value in the memory, and increasing the
				-- stack pointer for the address count.
				-----
				elsif currentState <= stateProcessLL then						-- Set the data and the address for storing the data to the output RAM.
					dataToSend <= inLL;
					addressToSend <= spLL;
					returnState <= stateProcessLLIncreaseSP;
				elsif currentState <= stateProcessLLIncreaseSP then		-- Increase the stack pointer for the LL component of the image
																							-- (raw data) which holds the approximation of the original image.
					spLL <= spLL + 1;
				
				
				
				-----
				-- Process the LH component of the image. This consists in counting the successive LH values which are lower than the given
				-- threshold, until a value that is >= THRESHOLD arrives.
				-----
				elsif currentState = stateProcessLHCount then				-- Increase the count of LH decomposed values which are lower than
																							-- the given threshold.
					sameCountLH <= sameCountLH + 1;
				elsif currentState = stateProcessLHSend1 then				-- Send the count of values which are lower than the threshold to
																							-- a location in the output RAM pointed to by the spLH stack pointer.
					if (inLH < THRESHOLD) then										-- If this condition is true, that means that sameCountLH is equal to
																							-- 255 and we jumped into this state because of the overflow, and not
																							-- because there was a valid data byte (inLH is not >= THRESHOLD).
																							-- We need to subtract 1 from the count, because we send the count
																							-- of zeros followed by a zero.
						dataToSend <= conv_std_logic_vector((sameCountLH - 1), (DATA_WIDTH));
					else
						dataToSend <= conv_std_logic_vector(sameCountLH, (DATA_WIDTH));
					end if;
					addressToSend <= spLH;
					returnState <= stateProcessLHIncreaseSP1;
				elsif currentState = stateProcessLHIncreaseSP1 then		-- Increase the LH stack pointer.
					spLH <= spLH + 1;
				elsif currentState = stateProcessLHSend2 then				-- Send the valid data byte that followed the sameCountLH (count of
																							-- values lower than the given threshold), or send a 0 if there was
																							-- an overflow in the count.
					if inLH < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inLH;
					end if;
					addressToSend <= spLH;
					returnState <= stateProcessLHIncreaseSP2;
				elsif currentState = stateProcessLHIncreaseSP2 then		-- Increase the LH stack pointer.
					spLH <= spLH + 1;
				elsif currentState = stateProcessLHClearCount then			-- Clear the count of values lower than the given threshold.
					sameCountLH <= 0;
					
				-----
				-- Process the HL component of the image (analogous to the LH component).
				-----
				elsif currentState = stateProcessHLCount then
					sameCountHL <= sameCountHL + 1;
				elsif currentState = stateProcessHLSend1 then
					if (inHL < THRESHOLD) then
						dataToSend <= conv_std_logic_vector((sameCountHL - 1), (DATA_WIDTH));
					else
						dataToSend <= conv_std_logic_vector(sameCountHL, (DATA_WIDTH));
					end if;
					addressToSend <= spHL;
					returnState <= stateProcessHLIncreaseSP1;
				elsif currentState = stateProcessHLIncreaseSP1 then
					spHL <= spHL + 1;
				elsif currentState = stateProcessHLSend2 then
					if inHL < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inHL;
					end if;
					addressToSend <= spHL;
					returnState <= stateProcessHLIncreaseSP2;
				elsif currentState = stateProcessHLIncreaseSP2 then
					spHL <= spHL + 1;
				elsif currentState = stateProcessHLClearCount then
					sameCountHL <= 0;

				-----
				-- Process the HH component of the image (analogous to the LH component).
				-----
				elsif currentState = stateProcessHHCount then
					sameCountHH <= sameCountHH + 1;
				elsif currentState = stateProcessHHSend1 then
					if (inHH < THRESHOLD) then
						dataToSend <= conv_std_logic_vector((sameCountHH - 1), (DATA_WIDTH));
					else
						dataToSend <= conv_std_logic_vector(sameCountHH, (DATA_WIDTH));
					end if;
					addressToSend <= spHH;
					returnState <= stateProcessHHIncreaseSP1;
				elsif currentState = stateProcessHHIncreaseSP1 then
					spHH <= spHH + 1;
				elsif currentState = stateProcessHHSend2 then
					if inHH < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inHH;
					end if;
					addressToSend <= spHH;
					returnState <= stateProcessHHIncreaseSP2;
				elsif currentState = stateProcessHHIncreaseSP2 then
					spHH <= spHH + 1;
				elsif currentState = stateProcessHHClearCount then
					sameCountHH <= 0;
				
					
				

				-----------------------------------------------------------------
				-- This section checks if there were trailing zeros
				-- at the end of the decomposition. In case that the
				-- last pixel was lesser than the threshold (which is
				-- very likely), the sameCount of a particular component
				-- would be higher than zero, and needs to be written
				-- after the control unit has finished decomposing the
				-- input image). These states execute only after the
				-- cuFinishedProcessing signal is set high.
				-----------------------------------------------------------------
				-----
				-- Process the LH component of the image.
				-----
				elsif currentState = stateSendRemainingDataLH1 then
					dataToSend <= conv_std_logic_vector(sameCountLH - 1, (DATA_WIDTH));
					addressToSend <= spLH;
					returnState <= stateSendRemainingDataLHIncreaseSP1;
				elsif currentState = stateSendRemainingDataLHIncreaseSP1 then
					spLH <= spLH + 1;
				elsif currentState = stateSendRemainingDataLH2 then
					if inLH < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inLH;
					end if;
					addressToSend <= spLH;
					returnState <= stateSendRemainingDataLHIncreaseSP2;
				elsif currentState = stateSendRemainingDataLHIncreaseSP2 then
					spLH <= spLH + 1;
				elsif currentState = stateSendRemainingDataLHClearCount then
					sameCountLH <= 0;

				-----
				-- Process the HL component of the image (same as LH).
				-----
				elsif currentState = stateSendRemainingDataHL1 then
					dataToSend <= conv_std_logic_vector(sameCountHL - 1, (DATA_WIDTH));
					addressToSend <= spHL;
					returnState <= stateSendRemainingDataHLIncreaseSP1;
				elsif currentState = stateSendRemainingDataHLIncreaseSP1 then
					spHL <= spHL + 1;
				elsif currentState = stateSendRemainingDataHL2 then
					if inHL < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inHL;
					end if;
					addressToSend <= spHL;
					returnState <= stateSendRemainingDataHLIncreaseSP2;
				elsif currentState = stateSendRemainingDataHLIncreaseSP2 then
					spHL <= spHL + 1;
				elsif currentState = stateSendRemainingDataHLClearCount then
					sameCountHL <= 0;
				
				-----
				-- Process the HH component of the image (same as LH).
				-----
				elsif currentState = stateSendRemainingDataHH1 then
					dataToSend <= conv_std_logic_vector(sameCountHH - 1, (DATA_WIDTH));
					addressToSend <= spHH;
					returnState <= stateSendRemainingDataHHIncreaseSP1;
				elsif currentState = stateSendRemainingDataHHIncreaseSP1 then
					spHH <= spHH + 1;
				elsif currentState = stateSendRemainingDataHH2 then
					if inHH < THRESHOLD then
						dataToSend <= (others => '0');
					else
						dataToSend <= inHH;
					end if;
					addressToSend <= spHH;
					returnState <= stateSendRemainingDataHHIncreaseSP2;
				elsif currentState = stateSendRemainingDataHHIncreaseSP2 then
					spHH <= spHH + 1;
				elsif currentState = stateSendRemainingDataHHClearCount then
					sameCountHH <= 0;
					
				
				-----------------------------------------------------------------
				-- After the image has been compressed, we need to move the
				-- HL and HH chunks right after the LH chunk, to make data
				-- contiguous. This is because between each of these components
				-- there is most likely a large number of zeros (which we need
				-- to remove in order to actually achieve compression).
				-----------------------------------------------------------------
				-----
				-- Move the HL component of the image
				-----
				elsif currentState = stateMoveHLReadData then
					dataToSend <= dataIn;
					addressToSend <= spLH;
					returnState <= stateMoveHLIncreaseSP;
				elsif currentState = stateMoveHLIncreaseSP then
					spHLMoving <= spHLMoving + 1;
					spLH <= spLH + 1;

				-----
				-- Move the HH component of the image (same as HL).
				-----
				elsif currentState = stateMoveHHReadData then
					dataToSend <= dataIn;
					addressToSend <= spLH;
					returnState <= stateMoveHHIncreaseSP;
				elsif currentState = stateMoveHHIncreaseSP then
					spHHMoving <= spHHMoving + 1;
					spLH <= spLH + 1;
					
					
					
				end if;
				
				currentState <= nextState;
			end if;
		end if;
	end process;
	
	-- Combinational part of the state machine.
	process (currentState, columnReady, rowReady, inLH, sameCountLH, inHL, sameCountHL, inHH, sameCountHH, addressToSend, dataToSend, returnState, cuFinishedProcessing, spHLMoving, spHHMoving, spLH, spHL, spHH)
	begin
		-- Set the default values for the signals in order to avoid generating latches.
		nextState <= stateReset;

		readyForNextData <= '0';
		address <= (others => '0');
		dataOut <= (others => '0');
		weOut <= '0';
		finishedCompressing <= '0';
		compressedDataSize <= (others => '0');

		case currentState is
			when stateReset =>											-- Initialize the state machine.
				nextState <= stateWaitForRowAndColumn;
			
			when stateWaitForRowAndColumn =>							-- Wait until the row and column ready signals are high.
																				-- These signals are used to decimate the output data.
																				-- Until both of these are high, we just loop through this state.
				readyForNextData <= '1';
				if ((rowReady = '1' and columnReady = '1') and cuFinishedProcessing = '0') then
					nextState <= stateProcessData;
				elsif (cuFinishedProcessing = '1') then
					nextState <= stateSendRemainingData;
				else
					nextState <= stateWaitForRowAndColumn;
				end if;
			
			
			
			-----------------------------------------------------------------
			-- These states are used for counting the values that are
			-- lower than the given threshold, and storing the results
			-- to the output RAM. These states occur while
			-- cuFinishedProcessing is low.
			-----------------------------------------------------------------
			-----
			-- Start processing the data.
			-----
			when stateProcessData =>
				nextState <= stateProcessLL;
				
			-----
			-- Process the LL component of the image. This consists simply of storing the raw value in the memory, and increasing the
			-- stack pointer for the address count.
			-----				
			when stateProcessLL =>
				nextState <= stateSendData;
			when stateProcessLLIncreaseSP =>
				nextState <= stateProcessLH;
				
			-----
			-- Process the LH component of the image. This consists in counting the successive LH values which are lower than the given
			-- threshold, until a value that is >= THRESHOLD arrives.
			-----					
			when stateProcessLH =>											-- Chech if the data value is lower than the given threshold, and
																					-- jump to appropriate states.
				if (inLH < conv_std_logic_vector(THRESHOLD, DATA_WIDTH)) then
					nextState <= stateProcessLHCount;
				else
					nextState <= stateProcessLHSend1;
				end if;
			when stateProcessLHCount =>									-- If the data value is lower than the threshold, increase the count.
				-- (In the synchronous process): Same count needs to be increased
				if (sameCountLH = 254) then								-- Check if the count will overflow. We compare with 254, because the
																					-- the count will be increased right before the state changes, from the
																					-- synchronous process of the state machine.
					nextState <= stateProcessLHSend1;
				else
					nextState <= stateProcessHL;
				end if;
			when stateProcessLHSend1 =>
				-- Here, the count of zeros (data lesser than threshold) is sent to RAM. Return state is set in the synchronous process (stateProcessLHIncreaseSP1).
				nextState <= stateSendData;
			when stateProcessLHIncreaseSP1 =>							-- Increase the stack pointer after storing the count.
				nextState <= stateProcessLHSend2;
			when stateProcessLHSend2 =>
				-- Here, the following data is sent to RAM. Return state is set in the synchronous process (stateProcessLHIncreaseSP2);
				nextState <= stateSendData;
			when stateProcessLHIncreaseSP2 =>							-- Increase the stack pointer after storing the data value.
				nextState <= stateProcessLHClearCount;
			when stateProcessLHClearCount =>								-- Clear the count, so it will be ready for the next batch of values.
				nextState <= stateProcessHL;
				
			-----
			-- Process the HL component of the image (analogous to the LH component).
			-----
			when stateProcessHL =>
				if (inHL <= conv_std_logic_vector(THRESHOLD, DATA_WIDTH)) then
					nextState <= stateProcessHLCount;
				else
					nextState <= stateProcessHLSend1;
				end if;
			when stateProcessHLCount =>
				-- (In the synchronous process): Same count needs to be increased
				if (sameCountHL = 254) then
					nextState <= stateProcessHLSend1;
				else
					nextState <= stateProcessHH;
				end if;
			when stateProcessHLSend1 =>
				-- Here, the count of zeros (data lesser than threshold) is sent to RAM. Return state is set in the synchronous process (stateProcessHLIncreaseSP1).
				nextState <= stateSendData;
			when stateProcessHLIncreaseSP1 =>
				nextState <= stateProcessHLSend2;
			when stateProcessHLSend2 =>
				-- Here, the following data is sent to RAM. Return state is set in the synchronous process (stateProcessHLIncreaseSP2);
				nextState <= stateSendData;
			when stateProcessHLIncreaseSP2 =>
				nextState <= stateProcessHLClearCount;
			when stateProcessHLClearCount =>
				nextState <= stateProcessHH;

			-----
			-- Process the HH component of the image (analogous to the LH component).
			-----
			when stateProcessHH =>
				if (inHH < conv_std_logic_vector(THRESHOLD, DATA_WIDTH)) then
					nextState <= stateProcessHHCount;
				else
					nextState <= stateProcessHHSend1;
				end if;
			when stateProcessHHCount =>
				-- (In the synchronous process): Same count needs to be increased
				if (sameCountHH = 254) then -- or cuFinishedProcessing = '1') then
					nextState <= stateProcessHHSend1;
				else
					nextState <= stateFinished;
				end if;
			when stateProcessHHSend1 =>
				-- Here, the count of zeros (data lesser than threshold) is sent to RAM. Return state is set in the synchronous process (stateProcessHHIncreaseSP1).
				nextState <= stateSendData;
			when stateProcessHHIncreaseSP1 =>
				nextState <= stateProcessHHSend2;
			when stateProcessHHSend2 =>
				-- Here, the following data is sent to RAM. Return state is set in the synchronous process (stateProcessHHIncreaseSP2);
				nextState <= stateSendData;
			when stateProcessHHIncreaseSP2 =>
				nextState <= stateProcessHHClearCount;
			when stateProcessHHClearCount =>
				nextState <= stateFinished;
			
			
			
			-----------------------------------------------------------------
			-- This section checks if there were trailing zeros
			-- at the end of the decomposition. In case that the
			-- last pixel was lesser than the threshold (which is
			-- very likely), the sameCount of a particular component
			-- would be higher than zero, and needs to be written
			-- after the control unit has finished decomposing the
			-- input image). These states execute only after the
			-- cuFinishedProcessing signal is set high.
			-----------------------------------------------------------------
			when stateSendRemainingData =>
				nextState <= stateSendRemainingDataLH1;
			
			-----
			-- Process the LH component of the image.
			-----
			when stateSendRemainingDataLH1 =>									-- Send the zero count if it exists, and jump
																							-- to stateSendRemainingDataLHIncreaseSP1 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataLHIncreaseSP1 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataLH2;
			when stateSendRemainingDataLH2 =>									-- Send the 0 data value, and jump
																							-- to stateSendRemainingDataLHIncreaseSP2 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataLHIncreaseSP2 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataLHClearCount;
			when stateSendRemainingDataLHClearCount =>						-- Be prudent, and clear the zero count.
				nextState <= stateSendRemainingDataHL1;

			-----
			-- Process the HL component of the image (same as LH).
			-----
			when stateSendRemainingDataHL1 =>									-- Send the zero count if it exists, and jump
																							-- to stateSendRemainingDataHLIncreaseSP1 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataHLIncreaseSP1 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataHL2;
			when stateSendRemainingDataHL2 =>									-- Send the 0 data value, and jump
																							-- to stateSendRemainingDataHLIncreaseSP2 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataHLIncreaseSP2 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataHLClearCount;
			when stateSendRemainingDataHLClearCount =>						-- Be prudent, and clear the zero count.
				nextState <= stateSendRemainingDataHH1;

			-----
			-- Process the HH component of the image (same as LH).
			-----
			when stateSendRemainingDataHH1 =>									-- Send the zero count if it exists, and jump
																							-- to stateSendRemainingDataHHIncreaseSP1 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataHHIncreaseSP1 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataHH2;
			when stateSendRemainingDataHH2 =>									-- Send the 0 data value, and jump
																							-- to stateSendRemainingDataHHIncreaseSP2 state afterwards
				nextState <= stateSendData;
			when stateSendRemainingDataHHIncreaseSP2 =>						-- Increase the stack pointer.
				nextState <= stateSendRemainingDataHHClearCount;
			when stateSendRemainingDataHHClearCount =>						-- Be prudent, and clear the zero count.
				nextState <= stateMoveHL;
			
			
			-----------------------------------------------------------------
			-- After the image has been compressed, we need to move the
			-- HL and HH chunks right after the LH chunk, to make data
			-- contiguous. This is because between each of these components
			-- there is most likely a large number of zeros (which we need
			-- to remove in order to actually achieve compression).
			-----------------------------------------------------------------
			-----
			-- Move the HL component of the image
			-----
			when stateMoveHL =>														-- Start moving the HL component of the image.
				nextState <= stateMoveHLCheckDone;
			when stateMoveHLCheckDone =>											-- Check if all data bytes have been moved, if so
																							-- jump to move the HH component.
				if (spHLMoving = spHL) then
					nextState <= stateMoveHH;
				else
					nextState <= stateMoveHLSetAddressRead;
				end if;
			when stateMoveHLSetAddressRead =>									-- Data byte has to first be read from memory. Set the
																							-- address of the current data byte that is to be moved
																							-- so we can read the contents at that address.
				address <= spHLMoving;
				nextState <= stateMoveHLReadData;
			when stateMoveHLReadData =>											-- Store the data byte to a register, and store it to the new location.
				nextState <= stateSendData;
			when stateMoveHLIncreaseSP =>											-- Increase the stack pointer pointing to the current contiguous
																							-- chunk of data (followed right after the LH component). Repeat
																							-- these states until all data bytes have been moved, then jump to
																							-- moving the HH component
				nextState <= stateMoveHLCheckDone;
			
			-----
			-- Move the HH component of the image (same as HL).
			-----
			when stateMoveHH =>														-- Start moving the HH component of the image.
				nextState <= stateMoveHHCheckDone;
			when stateMoveHHCheckDone =>											-- Check if all data bytes have been moved, if so
																							-- jump to the finished state.
				if (spHHMoving = spHH) then
					nextState <= stateFinished;
				else
					nextState <= stateMoveHHSetAddressRead;
				end if;
			when stateMoveHHSetAddressRead =>									-- Data byte has to first be read from memory. Set the
																							-- address of the current data byte that is to be moved
																							-- so we can read the contents at that address.
				address <= spHHMoving;
				nextState <= stateMoveHHReadData;
			when stateMoveHHReadData =>											-- Store the data byte to a register, and store it to the new location.
				nextState <= stateSendData;
			when stateMoveHHIncreaseSP =>											-- Increase the stack pointer pointing to the current contiguous
																							-- chunk of data (followed right after the LH component). Repeat
																							-- these states until all data bytes have been moved, then jump to
																							-- moving the HH component
				nextState <= stateMoveHHCheckDone;
			
			
			
			-----------------------------------------------------------------
			-- These are two general-purpose states for storing data to RAM.
			-- This operation is performed many times in this state machine
			-- so these states are used as a subroutine. The returnState
			-- signal MUST be set in the synchronous process of the design,
			-- otherwise unpredicted behaviour will occur.
			-----------------------------------------------------------------
			when stateSendData =>										-- Sets the address and the data to the corresponding busses.
																				-- Also enables writing to the output RAM.
				address <= addressToSend;
				dataOut <= dataToSend;
				weOut <= '1';
				nextState <= stateSendData2;
			when stateSendData2 =>										-- Disables writing to the output RAM and returns to a given state.
				weOut <= '0';
				nextState <= returnState;
				

			
			-----------------------------------------------------------------
			-- States which denote one of two things: either the current
			-- pixel has been processed, or all pixels have been processed
			-- (including moving of HL and LH data in memory).
			-----------------------------------------------------------------
			when stateFinished =>										-- This state is jumped to whenever the current pixel was processed.
				readyForNextData <= '1';
				nextState <= stateFinished2;
			when stateFinished2 =>										-- This state is used only as a 'wait' function, to allow the control
																				-- unit to settle its control signals.
				readyForNextData <= '1';
				nextState <= stateFinished3;
			when stateFinished3 =>										-- Check if the Control Unit has finished processing the data, if true,
																				-- then there is nothing else to do here and loop through this state.
																				-- Otherwise jump to the waiting state.
				readyForNextData <= '1';
				if (cuFinishedProcessing = '0') then
					nextState <= stateWaitForRowAndColumn;
				else
					finishedCompressing <= '1';
					compressedDataSize <= spLH;
					nextState <= stateFinished3;
				end if;
			end case;
	end process;
	
end Behavioral;
